library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.common_pkg.all;
use work.arith_pkg.all;

entity cpu is
    port (
        clock_i : in std_logic;
        reset_i : in std_logic;

        memoryAddress_o     : out std_logic_vector(15 downto 0);
        memoryReadData_i    :  in std_logic_vector(7 downto 0);
        memoryWriteData_o   : out std_logic_vector(7 downto 0);
        memoryWriteEnable_o : out std_logic
    );
end entity cpu;

architecture behavioral of cpu is

    signal instType_s : instruction_type;
    signal destType_s  : destination_type;
    signal srcType_s   : source_type;

    ------------------------------
    -- 16 bit register definitions
    signal pc_r     : std_logic_vector(15 downto 0);
    signal pcNext_r : std_logic_vector(15 downto 0);

    ------------------------------
    -- 8 bit register definitions.
    type regbank_type is array(natural range <>) of std_logic_vector(7 downto 0);

    -- Constants to directly select a register.
    constant REG_B   : std_logic_vector(2 downto 0) := "000";
    constant REG_C   : std_logic_vector(2 downto 0) := "001";
    constant REG_D   : std_logic_vector(2 downto 0) := "010";
    constant REG_E   : std_logic_vector(2 downto 0) := "011";
    constant REG_H   : std_logic_vector(2 downto 0) := "100";
    constant REG_L   : std_logic_vector(2 downto 0) := "101";
    constant REG_F   : std_logic_vector(2 downto 0) := "110";
    constant REG_A   : std_logic_vector(2 downto 0) := "110";

    -- This stores all the registers.
    signal regbank_r    : regbank_type(0 to 7);

    -- This holds data of the currently selected source register for reading.
    signal regReadData_s : std_logic_vector(7 downto 0);

    -- This selects the destination register (when destType_s = DEST_REGISTER).
    signal regDest_s    : std_logic_vector(2 downto 0);
    -- This selects the destination register (when srcType_s = SRC_REGISTER).
    signal regSrc_s    : std_logic_vector(2 downto 0);

    -- The result of the current calculation, will be written to the
    -- destination bus.
    signal result_s  : std_logic_vector(7 downto 0);

    -- The opcode register stores the opcode, obviously.
    -- The opcodeImm register stores an intermediate operand, if required.
    -- The opcode registers are delayed by one cycle.
    signal opcode_r    : std_logic_vector(7 downto 0);
    signal opcodeImm_r : std_logic_vector(7 downto 0);

    -- The signal variants are always valid thanks to an additional mux.
    signal opcode_s    : std_logic_vector(7 downto 0);
    signal opcodeImm_s : std_logic_vector(7 downto 0);

    -- The control signals of the CPU.
    -- Fetch our opcode, e.g. put the PC on the address bus.
    signal ctrlFetchOp_s     : std_logic;
    -- Decode the opcode, e.g. read the opcode register from the address bus.
    signal ctrlDecodeOp_s    : std_logic;
    -- Fetch an immediate operand
    signal ctrlFetchOpImm_s  : std_logic;
    -- Decode an immediate operand
    signal ctrlDecodeOpImm_s : std_logic;
    -- Increment the program counter
    signal ctrlIncPc_s       : std_logic;
    -- Execute the opcode
    signal ctrlExecute_s     : std_logic;

    -- This signal goes high when the current decoded opcode requires an
    -- immediate operand. This signal is generated by the decoder.
    signal requireImm_s : std_logic;

    type state_type is (
        STATE_FETCH,
        STATE_DECODE,
        STATE_DECODE_IMM
    );
    signal state_r     : state_type;
    signal stateNext_r : state_type;

    ----
    -- The original CPU is a bit slow, so we have several cycles per
    -- instruction available.
    -- Depending on the opcode, we have either 4, 8, 12 or 16 cycles available.
    -- The first two cycles are always the same:
    -- Stage 0: fetch the opcode by putting the program counter on the address
    --          bus. we also increment the program counter in this stage.
    -- Stage 1: the operand should now be on the data read bus, so we can
    --          decode it.
    -- Stage 2: here things get different depending on the opcode.
    --          * if the opcode requires an operand, we fetch it here.
    --          * otherwise we execute the opcode.
    -- Stage 3: if the opcode required an immidiate, it is executed here
    --          instead. Otherwise this stage is skipped.

begin

    -- The decoder instance. This component takes our opcode, decodes it and
    -- generates signals related to fetching more words.
    -- It generates a signal if we require an additional immediate value
    -- and if the opcode is complete or not.
    -- When the opcode is reported as completed, the type, source and
    -- destination signals can be used to execute the instruction.
    decoder_inst: entity work.decoder
        port map (
            clock_i       => clock_i,
            reset_i       => reset_i,

            -- The opcode we're decoding
            opcode_i      => opcode_s,

            -- When ready_o is high, this indicates the kind of instruction
            instType_o    => instType_s,
            srcType_o     => srcType_s,
            destType_o    => destType_s,

            -- The source and destination register indexes
            regDest_o     => regDest_s,
            regSrc_o      => regSrc_s,

            -- Inform the decoder that the opcode or immediate fields are read
            -- succesfully.
            opReady_i     => ctrlDecodeOp_s,
            immReady_i    => ctrlDecodeOpImm_s,

            ready_o       => ctrlExecute_s
        );

    -- The requested memory address. For now only the program counter is used
    -- when we fetch an opcode or an immediate.
    memoryAddress_o <= pc_r when ctrlFetchOp_s = '1' or ctrlFetchOpImm_s = '1'
                   else (others => 'Z');

    -- Writing is not done yet.
    memoryWriteEnable_o <= '0';

    -- Read the selected register.
    regReadData_s <= regbank_r(to_integer(unsigned(regSrc_s)));

    -- The result of our current operation, which will be written back.
    result_s <= opcodeImm_s   when srcType_s = SRC_IMMEDIATE
           else regReadData_s when srcType_s = SRC_REGISTER 
           else (others => '0');

    -- Bypass the opcode register when it is being decoded.
    opcode_s    <= memoryReadData_i when ctrlDecodeOp_s = '1'    else opcode_r;
    opcodeImm_s <= memoryReadData_i when ctrlDecodeOpImm_s = '1' else opcodeImm_r;

    -- The general clocked process, does state transitions and program counter
    -- incrementing.
    clock_proc: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            state_r <= STATE_FETCH;
            pc_r <= (others => '0');
        elsif rising_edge(clock_i) then
            pc_r <= pcNext_r;
            state_r <= stateNext_r;
        end if;
    end process;

    -- The register bank clocked process.
    reg_proc: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            regbank_r <= (others => (others => '0'));
        elsif rising_edge(clock_i) then
            if ctrlExecute_s = '1' and destType_s = DEST_REGISTER then
                regbank_r(to_integer(unsigned(regDest_s))) <= result_s;
            end if;
        end if;
    end process;

    -- The combinatorial state machine process.
    -- This produces the real control signals and calculates the next state,
    -- depending on the current state and if require an additional intermediate
    -- or not.
    state_comb_proc: process (state_r, srcType_s)
    begin
        stateNext_r <= state_r;
        ctrlFetchOp_s     <= '0';
        ctrlFetchOpImm_s  <= '0';
        ctrlDecodeOp_s    <= '0';
        ctrlDecodeOpImm_s <= '0';
        ctrlIncPc_s       <= '0';

        case state_r is
            -- The first stage fetches the opcode and increments the program
            -- counter.
            when STATE_FETCH  =>
                ctrlFetchOp_s <= '1';
                ctrlIncPc_s   <= '1';
                stateNext_r   <= STATE_DECODE;

            -- In the second state, the opcode is available and can be decoded.
            -- The decoder starts and notifies us if we require to fetch an
            -- additional byte.
            when STATE_DECODE =>
                -- Inform the decoder that the instruction is available.
                ctrlDecodeOp_s <= '1';

                -- Check if the decoder requires an additional intermediate.
                if srcType_s = SRC_IMMEDIATE then
                    -- Issue a fetch and increment of the program counter.
                    ctrlFetchOpImm_s <= '1';
                    ctrlIncPc_s <= '1';
                    stateNext_r <= STATE_DECODE_IMM;
                else
                    stateNext_r <= STATE_FETCH;
                end if;
            when STATE_DECODE_IMM =>
                -- Inform the decoder that the intermediate is available.
                ctrlDecodeOpImm_s <= '1';

                stateNext_r <= STATE_FETCH;

        end case;
    end process;

    -- This process stores the opcode or immediate values in their respective
    -- registers.
    opcode_reg_proc_s: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            opcode_r <= (others => '0');
        elsif rising_edge(clock_i) then
            if ctrlDecodeOp_s = '1' then
                opcode_r <= memoryReadData_i;
            end if;
            if ctrlDecodeOpImm_s = '1' then
                opcodeImm_r <= memoryReadData_i;
            end if;
        end if;
    end process;

    -- Calculate the next program counter.
    pc_next_proc: process (ctrlIncPc_s, pc_r)
    begin
        pcNext_r <= pc_r;
        if ctrlIncPc_s = '1' then
            pcNext_r <= increment(pc_r);
        end if;
    end process;

end architecture behavioral;
