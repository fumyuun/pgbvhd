library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cpu is
    port (
        clock_i : in std_logic;
        reset_i : in std_logic;

        memoryAddress_o     : out std_logic_vector(15 downto 0);
        memoryReadData_i    :  in std_logic_vector(7 downto 0);
        memoryWriteData_o   : out std_logic_vector(7 downto 0);
        memoryWriteEnable_o : out std_logic
    );
end entity cpu;

architecture behavioral of cpu is

    ------------------------------
    -- 16 bit register definitions
    signal pc_r     : std_logic_vector(15 downto 0);
    signal pcNext_r : std_logic_vector(15 downto 0);

    ------------------------------
    -- 8 bit register definitions.
    type regbank_type is array(natural range <>) of std_logic_vector(7 downto 0);

    -- Constants to directly select a register.
    constant REG_B   : std_logic_vector(2 downto 0) := "000";
    constant REG_C   : std_logic_vector(2 downto 0) := "001";
    constant REG_D   : std_logic_vector(2 downto 0) := "010";
    constant REG_E   : std_logic_vector(2 downto 0) := "011";
    constant REG_H   : std_logic_vector(2 downto 0) := "100";
    constant REG_L   : std_logic_vector(2 downto 0) := "101";
    constant REG_F   : std_logic_vector(2 downto 0) := "110";
    constant REG_A   : std_logic_vector(2 downto 0) := "110";

    -- This stores all the registers.
    signal regbank_r    : regbank_type(0 to 7);

    -- This selects the destination register.
    signal regDest_s    : std_logic_vector(2 downto 0);

    -- Write enable to the destination register.
    signal regWe_s      : std_logic;

    -- The result of the current calculation, will be written to the
    -- destination bus.
    signal result_s  : std_logic_vector(7 downto 0);

    -- The opcode register stores the opcode, obviously.
    -- The opcodeImm register stores an intermediate operand, if required.
    -- The opcode registers are delayed by one cycle.
    signal opcode_r    : std_logic_vector(7 downto 0);
    signal opcodeImm_r : std_logic_vector(7 downto 0);

    -- The signal variants are always valid thanks to an additional mux.
    signal opcode_s    : std_logic_vector(7 downto 0);
    signal opcodeImm_s : std_logic_vector(7 downto 0);

    -- The control signals of the CPU.
    -- Fetch our opcode, e.g. put the PC on the address bus.
    signal ctrlFetchOp_s     : std_logic;
    -- Decode the opcode, e.g. read the opcode register from the address bus.
    signal ctrlDecodeOp_s    : std_logic;
    -- Fetch an immediate operand
    signal ctrlFetchOpImm_s  : std_logic;
    -- Decode an immediate operand
    signal ctrlDecodeOpImm_s : std_logic;
    -- Increment the program counter
    signal ctrlIncPc_s       : std_logic;
    -- Execute the opcode
    signal ctrlExecute_s     : std_logic;

    -- This signal goes high when the current decoded opcode requires an
    -- immediate operand. This signal is generated by the decoder.
    signal requireImm_s : std_logic;

    type state_type is (
        STATE_FETCH,
        STATE_DECODE,
        STATE_DECODE_IMM
    );
    signal state_r     : state_type;
    signal stateNext_r : state_type;

    ----
    -- The original CPU is a bit slow, so we have several cycles per
    -- instruction available.
    -- Depending on the opcode, we have either 4, 8, 12 or 16 cycles available.
    -- The first two cycles are always the same:
    -- Stage 0: fetch the opcode by putting the program counter on the address
    --          bus. we also increment the program counter in this stage.
    -- Stage 1: the operand should now be on the data read bus, so we can
    --          decode it.
    -- Stage 2: here things get different depending on the opcode.
    --          * if the opcode requires an operand, we fetch it here.
    --          * otherwise we execute the opcode.
    -- Stage 3: if the opcode required an immidiate, it is executed here
    --          instead. Otherwise this stage is skipped.

begin

    decoder_inst: entity work.decoder
        port map (
            clock_i       => clock_i,
            reset_i       => reset_i,

            opcode_i      => opcode_s,

            regDest_o     => regDest_s,
            regWe_o       => regWe_s,

            opReady_i     => ctrlDecodeOp_s,
            immReady_i    => ctrlDecodeOpImm_s,

            requiresImm_o => requireImm_s,
            ready_o       => ctrlExecute_s
        );

    memoryAddress_o <= pc_r when ctrlFetchOp_s = '1' or ctrlFetchOpImm_s = '1'
                   else (others => 'Z');

    memoryWriteEnable_o <= '0';

    result_s <= opcodeImm_s when requireImm_s = '1' else (others => '0');

    -- Bypass the opcode register when it is being decoded.
    opcode_s     <= memoryReadData_i when ctrlDecodeOp_s = '1'     else opcode_r;
    opcodeImm_s <= memoryReadData_i when ctrlDecodeOpImm_s = '1' else opcodeImm_r;

    pc_reg_proc: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            pc_r <= (others => '0');
        elsif rising_edge(clock_i) then
            pc_r <= pcNext_r;
        end if;
    end process;

    reg_proc: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            regbank_r <= (others => (others => '0'));
        elsif rising_edge(clock_i) then
            if ctrlExecute_s = '1' and regWe_s = '1' then
                regbank_r(to_integer(unsigned(regDest_s))) <= result_s;
            end if;
        end if;
    end process;

    state_reg_proc: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            state_r <= STATE_FETCH;
        elsif rising_edge(clock_i) then
            state_r <= stateNext_r;
        end if;
    end process;

    state_comb_proc: process (state_r, requireImm_s)
    begin
        stateNext_r <= state_r;
        ctrlFetchOp_s      <= '0';
        ctrlFetchOpImm_s  <= '0';
        ctrlDecodeOp_s     <= '0';
        ctrlDecodeOpImm_s <= '0';
        ctrlIncPc_s        <= '0';

        case state_r is
            when STATE_FETCH  =>
                ctrlFetchOp_s <= '1';
                ctrlIncPc_s    <= '1';
                stateNext_r <= STATE_DECODE;

            when STATE_DECODE => 
                ctrlDecodeOp_s <= '1';

                if requireImm_s = '1' then
                    ctrlFetchOpImm_s <= '1';
                    ctrlIncPc_s <= '1';
                    stateNext_r <= STATE_DECODE_IMM;
                else
                    stateNext_r <= STATE_FETCH;
                end if;
            when STATE_DECODE_IMM =>
                ctrlDecodeOpImm_s <= '1';

                stateNext_r <= STATE_FETCH;

        end case;
    end process;

    opcode_reg_proc_s: process (reset_i, clock_i)
    begin
        if reset_i = '1' then
            opcode_r <= (others => '0');
        elsif rising_edge(clock_i) then
            if ctrlDecodeOp_s = '1' then
                opcode_r <= memoryReadData_i;
            end if;
            if ctrlDecodeOpImm_s = '1' then
                opcodeImm_r <= memoryReadData_i;
            end if;
        end if;
    end process;

    pc_next_proc: process (ctrlIncPc_s, pc_r)
    begin
        pcNext_r <= pc_r;
        if ctrlIncPc_s = '1' then
            pcNext_r <= std_logic_vector(to_unsigned(to_integer(unsigned(pc_r) + 1), pcNext_r'length));
        end if;
    end process;

end architecture behavioral;
